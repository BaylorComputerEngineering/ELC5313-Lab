`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/08/2025 02:58:22 PM
// Design Name: 
// Module Name: mod3counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mod3counter (
    input  logic [1:0] num,
    output logic [1:0] mod3num
);
    always_comb begin

    // TODO: implement modulo-3 logic
    
    end
endmodule
